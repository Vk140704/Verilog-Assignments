//13. Create a simple ALU module using only blocking assignments.
