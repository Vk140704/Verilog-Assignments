// /*10.Part Select Operation
// Extract lower nibble from reg [7:0] bus using bus[3:0].*/
// module part_select
//   reg [7:0]bus;
//   initial begin
//     data= 8'b00101010;
//     assign d= bus[3:0];
//   end 

// endmodule 

reg [7:0]bus;
int a;
initial begin
  if (bus[i]>4);
  a=0;
  else 
    a=a+1;
  
end
