	//1bit full adder
	module full_adder(
	 input a,b,cin,
       	 output sum,cout);
	wire g,x,y,z;

	xor(g,a,b);
	xor(sum,cin,g);
	and(x,a,b);
	and(y,b,cin);
	and(z,cin,a);
	or(cout,x,y,z);

   endmodule

   // 4-bit ripple carry adder
      module rca4bit(
	input [3:0]a,b,
	input cin,
	output [3:0]sum);
     wire c0,c1,c2;

full_adder fa0(.a(a[0]),.b(b[0]),.cin(cin[0]),,.sum(sum[0]),.cout(c0));
full_adder fa1(.a(a[1]),.b(b[1]),.cin(c0),.sum(sum[1]),.cout(c1));
full_adder fa2(.a(a[2]),.b(b[2]),.cin(c1),.sum(sum[2]),.cout(c2));
full_adder fa3(.a(a[3]),.b(b[3]),.cin(c2),.sum(sum[3]),.cout(cout));
endmodule
