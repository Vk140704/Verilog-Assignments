module nor_gate (input a,b,output f);
  nor(f,a,b);
endmodule
